module prog(adres,out);

input [4:0] adres;
output [31:0] out;
reg [31:0] out;
 
reg [31:0] pmem [31:0];

always @(*)

begin
	out=pmem[adres];
end

initial
begin
pmem[0]=32'b10000000010000000000000000000001;
pmem[1]=32'b10000000100000000000000000000010;
pmem[2]=32'b10000000110000000000000000000011;
pmem[3]=32'b10000001000000000000000000000100;
pmem[4]=32'b00110001010000000000000000100010;
pmem[5]=32'b00101001100000000000000010100011;
pmem[6]=32'b00110001110000000000000011000100;
end

endmodule